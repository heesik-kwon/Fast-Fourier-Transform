`timescale 1ns / 1ps

module twf_m0_rom (
    input  logic              clk,
    input  logic        [8:0] addr,
    output logic signed [9:0] w_re,
    output logic signed [9:0] w_im
);

    always_ff @(posedge clk) begin
        case (addr)
            9'd0: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd1: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd2: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd3: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd4: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd5: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd6: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd7: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd8: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd9: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd10: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd11: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd12: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd13: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd14: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd15: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd16: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd17: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd18: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd19: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd20: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd21: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd22: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd23: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd24: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd25: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd26: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd27: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd28: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd29: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd30: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd31: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd32: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd33: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd34: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd35: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd36: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd37: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd38: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd39: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd40: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd41: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd42: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd43: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd44: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd45: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd46: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd47: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd48: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd49: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd50: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd51: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd52: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd53: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd54: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd55: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd56: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd57: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd58: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd59: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd60: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd61: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd62: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd63: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd64: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd65: begin
                w_re = 10'sd128;
                w_im = -10'sd6;
            end
            9'd66: begin
                w_re = 10'sd127;
                w_im = -10'sd13;
            end
            9'd67: begin
                w_re = 10'sd127;
                w_im = -10'sd19;
            end
            9'd68: begin
                w_re = 10'sd126;
                w_im = -10'sd25;
            end
            9'd69: begin
                w_re = 10'sd124;
                w_im = -10'sd31;
            end
            9'd70: begin
                w_re = 10'sd122;
                w_im = -10'sd37;
            end
            9'd71: begin
                w_re = 10'sd121;
                w_im = -10'sd43;
            end
            9'd72: begin
                w_re = 10'sd118;
                w_im = -10'sd49;
            end
            9'd73: begin
                w_re = 10'sd116;
                w_im = -10'sd55;
            end
            9'd74: begin
                w_re = 10'sd113;
                w_im = -10'sd60;
            end
            9'd75: begin
                w_re = 10'sd110;
                w_im = -10'sd66;
            end
            9'd76: begin
                w_re = 10'sd106;
                w_im = -10'sd71;
            end
            9'd77: begin
                w_re = 10'sd103;
                w_im = -10'sd76;
            end
            9'd78: begin
                w_re = 10'sd99;
                w_im = -10'sd81;
            end
            9'd79: begin
                w_re = 10'sd95;
                w_im = -10'sd86;
            end
            9'd80: begin
                w_re = 10'sd91;
                w_im = -10'sd91;
            end
            9'd81: begin
                w_re = 10'sd86;
                w_im = -10'sd95;
            end
            9'd82: begin
                w_re = 10'sd81;
                w_im = -10'sd99;
            end
            9'd83: begin
                w_re = 10'sd76;
                w_im = -10'sd103;
            end
            9'd84: begin
                w_re = 10'sd71;
                w_im = -10'sd106;
            end
            9'd85: begin
                w_re = 10'sd66;
                w_im = -10'sd110;
            end
            9'd86: begin
                w_re = 10'sd60;
                w_im = -10'sd113;
            end
            9'd87: begin
                w_re = 10'sd55;
                w_im = -10'sd116;
            end
            9'd88: begin
                w_re = 10'sd49;
                w_im = -10'sd118;
            end
            9'd89: begin
                w_re = 10'sd43;
                w_im = -10'sd121;
            end
            9'd90: begin
                w_re = 10'sd37;
                w_im = -10'sd122;
            end
            9'd91: begin
                w_re = 10'sd31;
                w_im = -10'sd124;
            end
            9'd92: begin
                w_re = 10'sd25;
                w_im = -10'sd126;
            end
            9'd93: begin
                w_re = 10'sd19;
                w_im = -10'sd127;
            end
            9'd94: begin
                w_re = 10'sd13;
                w_im = -10'sd127;
            end
            9'd95: begin
                w_re = 10'sd6;
                w_im = -10'sd128;
            end
            9'd96: begin
                w_re = 10'sd0;
                w_im = -10'sd128;
            end
            9'd97: begin
                w_re = -10'sd6;
                w_im = -10'sd128;
            end
            9'd98: begin
                w_re = -10'sd13;
                w_im = -10'sd127;
            end
            9'd99: begin
                w_re = -10'sd19;
                w_im = -10'sd127;
            end
            9'd100: begin
                w_re = -10'sd25;
                w_im = -10'sd126;
            end
            9'd101: begin
                w_re = -10'sd31;
                w_im = -10'sd124;
            end
            9'd102: begin
                w_re = -10'sd37;
                w_im = -10'sd122;
            end
            9'd103: begin
                w_re = -10'sd43;
                w_im = -10'sd121;
            end
            9'd104: begin
                w_re = -10'sd49;
                w_im = -10'sd118;
            end
            9'd105: begin
                w_re = -10'sd55;
                w_im = -10'sd116;
            end
            9'd106: begin
                w_re = -10'sd60;
                w_im = -10'sd113;
            end
            9'd107: begin
                w_re = -10'sd66;
                w_im = -10'sd110;
            end
            9'd108: begin
                w_re = -10'sd71;
                w_im = -10'sd106;
            end
            9'd109: begin
                w_re = -10'sd76;
                w_im = -10'sd103;
            end
            9'd110: begin
                w_re = -10'sd81;
                w_im = -10'sd99;
            end
            9'd111: begin
                w_re = -10'sd86;
                w_im = -10'sd95;
            end
            9'd112: begin
                w_re = -10'sd91;
                w_im = -10'sd91;
            end
            9'd113: begin
                w_re = -10'sd95;
                w_im = -10'sd86;
            end
            9'd114: begin
                w_re = -10'sd99;
                w_im = -10'sd81;
            end
            9'd115: begin
                w_re = -10'sd103;
                w_im = -10'sd76;
            end
            9'd116: begin
                w_re = -10'sd106;
                w_im = -10'sd71;
            end
            9'd117: begin
                w_re = -10'sd110;
                w_im = -10'sd66;
            end
            9'd118: begin
                w_re = -10'sd113;
                w_im = -10'sd60;
            end
            9'd119: begin
                w_re = -10'sd116;
                w_im = -10'sd55;
            end
            9'd120: begin
                w_re = -10'sd118;
                w_im = -10'sd49;
            end
            9'd121: begin
                w_re = -10'sd121;
                w_im = -10'sd43;
            end
            9'd122: begin
                w_re = -10'sd122;
                w_im = -10'sd37;
            end
            9'd123: begin
                w_re = -10'sd124;
                w_im = -10'sd31;
            end
            9'd124: begin
                w_re = -10'sd126;
                w_im = -10'sd25;
            end
            9'd125: begin
                w_re = -10'sd127;
                w_im = -10'sd19;
            end
            9'd126: begin
                w_re = -10'sd127;
                w_im = -10'sd13;
            end
            9'd127: begin
                w_re = -10'sd128;
                w_im = -10'sd6;
            end
            9'd128: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd129: begin
                w_re = 10'sd128;
                w_im = -10'sd3;
            end
            9'd130: begin
                w_re = 10'sd128;
                w_im = -10'sd6;
            end
            9'd131: begin
                w_re = 10'sd128;
                w_im = -10'sd9;
            end
            9'd132: begin
                w_re = 10'sd127;
                w_im = -10'sd13;
            end
            9'd133: begin
                w_re = 10'sd127;
                w_im = -10'sd16;
            end
            9'd134: begin
                w_re = 10'sd127;
                w_im = -10'sd19;
            end
            9'd135: begin
                w_re = 10'sd126;
                w_im = -10'sd22;
            end
            9'd136: begin
                w_re = 10'sd126;
                w_im = -10'sd25;
            end
            9'd137: begin
                w_re = 10'sd125;
                w_im = -10'sd28;
            end
            9'd138: begin
                w_re = 10'sd124;
                w_im = -10'sd31;
            end
            9'd139: begin
                w_re = 10'sd123;
                w_im = -10'sd34;
            end
            9'd140: begin
                w_re = 10'sd122;
                w_im = -10'sd37;
            end
            9'd141: begin
                w_re = 10'sd122;
                w_im = -10'sd40;
            end
            9'd142: begin
                w_re = 10'sd121;
                w_im = -10'sd43;
            end
            9'd143: begin
                w_re = 10'sd119;
                w_im = -10'sd46;
            end
            9'd144: begin
                w_re = 10'sd118;
                w_im = -10'sd49;
            end
            9'd145: begin
                w_re = 10'sd117;
                w_im = -10'sd52;
            end
            9'd146: begin
                w_re = 10'sd116;
                w_im = -10'sd55;
            end
            9'd147: begin
                w_re = 10'sd114;
                w_im = -10'sd58;
            end
            9'd148: begin
                w_re = 10'sd113;
                w_im = -10'sd60;
            end
            9'd149: begin
                w_re = 10'sd111;
                w_im = -10'sd63;
            end
            9'd150: begin
                w_re = 10'sd110;
                w_im = -10'sd66;
            end
            9'd151: begin
                w_re = 10'sd108;
                w_im = -10'sd68;
            end
            9'd152: begin
                w_re = 10'sd106;
                w_im = -10'sd71;
            end
            9'd153: begin
                w_re = 10'sd105;
                w_im = -10'sd74;
            end
            9'd154: begin
                w_re = 10'sd103;
                w_im = -10'sd76;
            end
            9'd155: begin
                w_re = 10'sd101;
                w_im = -10'sd79;
            end
            9'd156: begin
                w_re = 10'sd99;
                w_im = -10'sd81;
            end
            9'd157: begin
                w_re = 10'sd97;
                w_im = -10'sd84;
            end
            9'd158: begin
                w_re = 10'sd95;
                w_im = -10'sd86;
            end
            9'd159: begin
                w_re = 10'sd93;
                w_im = -10'sd88;
            end
            9'd160: begin
                w_re = 10'sd91;
                w_im = -10'sd91;
            end
            9'd161: begin
                w_re = 10'sd88;
                w_im = -10'sd93;
            end
            9'd162: begin
                w_re = 10'sd86;
                w_im = -10'sd95;
            end
            9'd163: begin
                w_re = 10'sd84;
                w_im = -10'sd97;
            end
            9'd164: begin
                w_re = 10'sd81;
                w_im = -10'sd99;
            end
            9'd165: begin
                w_re = 10'sd79;
                w_im = -10'sd101;
            end
            9'd166: begin
                w_re = 10'sd76;
                w_im = -10'sd103;
            end
            9'd167: begin
                w_re = 10'sd74;
                w_im = -10'sd105;
            end
            9'd168: begin
                w_re = 10'sd71;
                w_im = -10'sd106;
            end
            9'd169: begin
                w_re = 10'sd68;
                w_im = -10'sd108;
            end
            9'd170: begin
                w_re = 10'sd66;
                w_im = -10'sd110;
            end
            9'd171: begin
                w_re = 10'sd63;
                w_im = -10'sd111;
            end
            9'd172: begin
                w_re = 10'sd60;
                w_im = -10'sd113;
            end
            9'd173: begin
                w_re = 10'sd58;
                w_im = -10'sd114;
            end
            9'd174: begin
                w_re = 10'sd55;
                w_im = -10'sd116;
            end
            9'd175: begin
                w_re = 10'sd52;
                w_im = -10'sd117;
            end
            9'd176: begin
                w_re = 10'sd49;
                w_im = -10'sd118;
            end
            9'd177: begin
                w_re = 10'sd46;
                w_im = -10'sd119;
            end
            9'd178: begin
                w_re = 10'sd43;
                w_im = -10'sd121;
            end
            9'd179: begin
                w_re = 10'sd40;
                w_im = -10'sd122;
            end
            9'd180: begin
                w_re = 10'sd37;
                w_im = -10'sd122;
            end
            9'd181: begin
                w_re = 10'sd34;
                w_im = -10'sd123;
            end
            9'd182: begin
                w_re = 10'sd31;
                w_im = -10'sd124;
            end
            9'd183: begin
                w_re = 10'sd28;
                w_im = -10'sd125;
            end
            9'd184: begin
                w_re = 10'sd25;
                w_im = -10'sd126;
            end
            9'd185: begin
                w_re = 10'sd22;
                w_im = -10'sd126;
            end
            9'd186: begin
                w_re = 10'sd19;
                w_im = -10'sd127;
            end
            9'd187: begin
                w_re = 10'sd16;
                w_im = -10'sd127;
            end
            9'd188: begin
                w_re = 10'sd13;
                w_im = -10'sd127;
            end
            9'd189: begin
                w_re = 10'sd9;
                w_im = -10'sd128;
            end
            9'd190: begin
                w_re = 10'sd6;
                w_im = -10'sd128;
            end
            9'd191: begin
                w_re = 10'sd3;
                w_im = -10'sd128;
            end
            9'd192: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd193: begin
                w_re = 10'sd128;
                w_im = -10'sd9;
            end
            9'd194: begin
                w_re = 10'sd127;
                w_im = -10'sd19;
            end
            9'd195: begin
                w_re = 10'sd125;
                w_im = -10'sd28;
            end
            9'd196: begin
                w_re = 10'sd122;
                w_im = -10'sd37;
            end
            9'd197: begin
                w_re = 10'sd119;
                w_im = -10'sd46;
            end
            9'd198: begin
                w_re = 10'sd116;
                w_im = -10'sd55;
            end
            9'd199: begin
                w_re = 10'sd111;
                w_im = -10'sd63;
            end
            9'd200: begin
                w_re = 10'sd106;
                w_im = -10'sd71;
            end
            9'd201: begin
                w_re = 10'sd101;
                w_im = -10'sd79;
            end
            9'd202: begin
                w_re = 10'sd95;
                w_im = -10'sd86;
            end
            9'd203: begin
                w_re = 10'sd88;
                w_im = -10'sd93;
            end
            9'd204: begin
                w_re = 10'sd81;
                w_im = -10'sd99;
            end
            9'd205: begin
                w_re = 10'sd74;
                w_im = -10'sd105;
            end
            9'd206: begin
                w_re = 10'sd66;
                w_im = -10'sd110;
            end
            9'd207: begin
                w_re = 10'sd58;
                w_im = -10'sd114;
            end
            9'd208: begin
                w_re = 10'sd49;
                w_im = -10'sd118;
            end
            9'd209: begin
                w_re = 10'sd40;
                w_im = -10'sd122;
            end
            9'd210: begin
                w_re = 10'sd31;
                w_im = -10'sd124;
            end
            9'd211: begin
                w_re = 10'sd22;
                w_im = -10'sd126;
            end
            9'd212: begin
                w_re = 10'sd13;
                w_im = -10'sd127;
            end
            9'd213: begin
                w_re = 10'sd3;
                w_im = -10'sd128;
            end
            9'd214: begin
                w_re = -10'sd6;
                w_im = -10'sd128;
            end
            9'd215: begin
                w_re = -10'sd16;
                w_im = -10'sd127;
            end
            9'd216: begin
                w_re = -10'sd25;
                w_im = -10'sd126;
            end
            9'd217: begin
                w_re = -10'sd34;
                w_im = -10'sd123;
            end
            9'd218: begin
                w_re = -10'sd43;
                w_im = -10'sd121;
            end
            9'd219: begin
                w_re = -10'sd52;
                w_im = -10'sd117;
            end
            9'd220: begin
                w_re = -10'sd60;
                w_im = -10'sd113;
            end
            9'd221: begin
                w_re = -10'sd68;
                w_im = -10'sd108;
            end
            9'd222: begin
                w_re = -10'sd76;
                w_im = -10'sd103;
            end
            9'd223: begin
                w_re = -10'sd84;
                w_im = -10'sd97;
            end
            9'd224: begin
                w_re = -10'sd91;
                w_im = -10'sd91;
            end
            9'd225: begin
                w_re = -10'sd97;
                w_im = -10'sd84;
            end
            9'd226: begin
                w_re = -10'sd103;
                w_im = -10'sd76;
            end
            9'd227: begin
                w_re = -10'sd108;
                w_im = -10'sd68;
            end
            9'd228: begin
                w_re = -10'sd113;
                w_im = -10'sd60;
            end
            9'd229: begin
                w_re = -10'sd117;
                w_im = -10'sd52;
            end
            9'd230: begin
                w_re = -10'sd121;
                w_im = -10'sd43;
            end
            9'd231: begin
                w_re = -10'sd123;
                w_im = -10'sd34;
            end
            9'd232: begin
                w_re = -10'sd126;
                w_im = -10'sd25;
            end
            9'd233: begin
                w_re = -10'sd127;
                w_im = -10'sd16;
            end
            9'd234: begin
                w_re = -10'sd128;
                w_im = -10'sd6;
            end
            9'd235: begin
                w_re = -10'sd128;
                w_im = 10'sd3;
            end
            9'd236: begin
                w_re = -10'sd127;
                w_im = 10'sd13;
            end
            9'd237: begin
                w_re = -10'sd126;
                w_im = 10'sd22;
            end
            9'd238: begin
                w_re = -10'sd124;
                w_im = 10'sd31;
            end
            9'd239: begin
                w_re = -10'sd122;
                w_im = 10'sd40;
            end
            9'd240: begin
                w_re = -10'sd118;
                w_im = 10'sd49;
            end
            9'd241: begin
                w_re = -10'sd114;
                w_im = 10'sd58;
            end
            9'd242: begin
                w_re = -10'sd110;
                w_im = 10'sd66;
            end
            9'd243: begin
                w_re = -10'sd105;
                w_im = 10'sd74;
            end
            9'd244: begin
                w_re = -10'sd99;
                w_im = 10'sd81;
            end
            9'd245: begin
                w_re = -10'sd93;
                w_im = 10'sd88;
            end
            9'd246: begin
                w_re = -10'sd86;
                w_im = 10'sd95;
            end
            9'd247: begin
                w_re = -10'sd79;
                w_im = 10'sd101;
            end
            9'd248: begin
                w_re = -10'sd71;
                w_im = 10'sd106;
            end
            9'd249: begin
                w_re = -10'sd63;
                w_im = 10'sd111;
            end
            9'd250: begin
                w_re = -10'sd55;
                w_im = 10'sd116;
            end
            9'd251: begin
                w_re = -10'sd46;
                w_im = 10'sd119;
            end
            9'd252: begin
                w_re = -10'sd37;
                w_im = 10'sd122;
            end
            9'd253: begin
                w_re = -10'sd28;
                w_im = 10'sd125;
            end
            9'd254: begin
                w_re = -10'sd19;
                w_im = 10'sd127;
            end
            9'd255: begin
                w_re = -10'sd9;
                w_im = 10'sd128;
            end
            9'd256: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd257: begin
                w_re = 10'sd128;
                w_im = -10'sd2;
            end
            9'd258: begin
                w_re = 10'sd128;
                w_im = -10'sd3;
            end
            9'd259: begin
                w_re = 10'sd128;
                w_im = -10'sd5;
            end
            9'd260: begin
                w_re = 10'sd128;
                w_im = -10'sd6;
            end
            9'd261: begin
                w_re = 10'sd128;
                w_im = -10'sd8;
            end
            9'd262: begin
                w_re = 10'sd128;
                w_im = -10'sd9;
            end
            9'd263: begin
                w_re = 10'sd128;
                w_im = -10'sd11;
            end
            9'd264: begin
                w_re = 10'sd127;
                w_im = -10'sd13;
            end
            9'd265: begin
                w_re = 10'sd127;
                w_im = -10'sd14;
            end
            9'd266: begin
                w_re = 10'sd127;
                w_im = -10'sd16;
            end
            9'd267: begin
                w_re = 10'sd127;
                w_im = -10'sd17;
            end
            9'd268: begin
                w_re = 10'sd127;
                w_im = -10'sd19;
            end
            9'd269: begin
                w_re = 10'sd126;
                w_im = -10'sd20;
            end
            9'd270: begin
                w_re = 10'sd126;
                w_im = -10'sd22;
            end
            9'd271: begin
                w_re = 10'sd126;
                w_im = -10'sd23;
            end
            9'd272: begin
                w_re = 10'sd126;
                w_im = -10'sd25;
            end
            9'd273: begin
                w_re = 10'sd125;
                w_im = -10'sd27;
            end
            9'd274: begin
                w_re = 10'sd125;
                w_im = -10'sd28;
            end
            9'd275: begin
                w_re = 10'sd125;
                w_im = -10'sd30;
            end
            9'd276: begin
                w_re = 10'sd124;
                w_im = -10'sd31;
            end
            9'd277: begin
                w_re = 10'sd124;
                w_im = -10'sd33;
            end
            9'd278: begin
                w_re = 10'sd123;
                w_im = -10'sd34;
            end
            9'd279: begin
                w_re = 10'sd123;
                w_im = -10'sd36;
            end
            9'd280: begin
                w_re = 10'sd122;
                w_im = -10'sd37;
            end
            9'd281: begin
                w_re = 10'sd122;
                w_im = -10'sd39;
            end
            9'd282: begin
                w_re = 10'sd122;
                w_im = -10'sd40;
            end
            9'd283: begin
                w_re = 10'sd121;
                w_im = -10'sd42;
            end
            9'd284: begin
                w_re = 10'sd121;
                w_im = -10'sd43;
            end
            9'd285: begin
                w_re = 10'sd120;
                w_im = -10'sd45;
            end
            9'd286: begin
                w_re = 10'sd119;
                w_im = -10'sd46;
            end
            9'd287: begin
                w_re = 10'sd119;
                w_im = -10'sd48;
            end
            9'd288: begin
                w_re = 10'sd118;
                w_im = -10'sd49;
            end
            9'd289: begin
                w_re = 10'sd118;
                w_im = -10'sd50;
            end
            9'd290: begin
                w_re = 10'sd117;
                w_im = -10'sd52;
            end
            9'd291: begin
                w_re = 10'sd116;
                w_im = -10'sd53;
            end
            9'd292: begin
                w_re = 10'sd116;
                w_im = -10'sd55;
            end
            9'd293: begin
                w_re = 10'sd115;
                w_im = -10'sd56;
            end
            9'd294: begin
                w_re = 10'sd114;
                w_im = -10'sd58;
            end
            9'd295: begin
                w_re = 10'sd114;
                w_im = -10'sd59;
            end
            9'd296: begin
                w_re = 10'sd113;
                w_im = -10'sd60;
            end
            9'd297: begin
                w_re = 10'sd112;
                w_im = -10'sd62;
            end
            9'd298: begin
                w_re = 10'sd111;
                w_im = -10'sd63;
            end
            9'd299: begin
                w_re = 10'sd111;
                w_im = -10'sd64;
            end
            9'd300: begin
                w_re = 10'sd110;
                w_im = -10'sd66;
            end
            9'd301: begin
                w_re = 10'sd109;
                w_im = -10'sd67;
            end
            9'd302: begin
                w_re = 10'sd108;
                w_im = -10'sd68;
            end
            9'd303: begin
                w_re = 10'sd107;
                w_im = -10'sd70;
            end
            9'd304: begin
                w_re = 10'sd106;
                w_im = -10'sd71;
            end
            9'd305: begin
                w_re = 10'sd106;
                w_im = -10'sd72;
            end
            9'd306: begin
                w_re = 10'sd105;
                w_im = -10'sd74;
            end
            9'd307: begin
                w_re = 10'sd104;
                w_im = -10'sd75;
            end
            9'd308: begin
                w_re = 10'sd103;
                w_im = -10'sd76;
            end
            9'd309: begin
                w_re = 10'sd102;
                w_im = -10'sd78;
            end
            9'd310: begin
                w_re = 10'sd101;
                w_im = -10'sd79;
            end
            9'd311: begin
                w_re = 10'sd100;
                w_im = -10'sd80;
            end
            9'd312: begin
                w_re = 10'sd99;
                w_im = -10'sd81;
            end
            9'd313: begin
                w_re = 10'sd98;
                w_im = -10'sd82;
            end
            9'd314: begin
                w_re = 10'sd97;
                w_im = -10'sd84;
            end
            9'd315: begin
                w_re = 10'sd96;
                w_im = -10'sd85;
            end
            9'd316: begin
                w_re = 10'sd95;
                w_im = -10'sd86;
            end
            9'd317: begin
                w_re = 10'sd94;
                w_im = -10'sd87;
            end
            9'd318: begin
                w_re = 10'sd93;
                w_im = -10'sd88;
            end
            9'd319: begin
                w_re = 10'sd92;
                w_im = -10'sd89;
            end
            9'd320: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd321: begin
                w_re = 10'sd128;
                w_im = -10'sd8;
            end
            9'd322: begin
                w_re = 10'sd127;
                w_im = -10'sd16;
            end
            9'd323: begin
                w_re = 10'sd126;
                w_im = -10'sd23;
            end
            9'd324: begin
                w_re = 10'sd124;
                w_im = -10'sd31;
            end
            9'd325: begin
                w_re = 10'sd122;
                w_im = -10'sd39;
            end
            9'd326: begin
                w_re = 10'sd119;
                w_im = -10'sd46;
            end
            9'd327: begin
                w_re = 10'sd116;
                w_im = -10'sd53;
            end
            9'd328: begin
                w_re = 10'sd113;
                w_im = -10'sd60;
            end
            9'd329: begin
                w_re = 10'sd109;
                w_im = -10'sd67;
            end
            9'd330: begin
                w_re = 10'sd105;
                w_im = -10'sd74;
            end
            9'd331: begin
                w_re = 10'sd100;
                w_im = -10'sd80;
            end
            9'd332: begin
                w_re = 10'sd95;
                w_im = -10'sd86;
            end
            9'd333: begin
                w_re = 10'sd89;
                w_im = -10'sd92;
            end
            9'd334: begin
                w_re = 10'sd84;
                w_im = -10'sd97;
            end
            9'd335: begin
                w_re = 10'sd78;
                w_im = -10'sd102;
            end
            9'd336: begin
                w_re = 10'sd71;
                w_im = -10'sd106;
            end
            9'd337: begin
                w_re = 10'sd64;
                w_im = -10'sd111;
            end
            9'd338: begin
                w_re = 10'sd58;
                w_im = -10'sd114;
            end
            9'd339: begin
                w_re = 10'sd50;
                w_im = -10'sd118;
            end
            9'd340: begin
                w_re = 10'sd43;
                w_im = -10'sd121;
            end
            9'd341: begin
                w_re = 10'sd36;
                w_im = -10'sd123;
            end
            9'd342: begin
                w_re = 10'sd28;
                w_im = -10'sd125;
            end
            9'd343: begin
                w_re = 10'sd20;
                w_im = -10'sd126;
            end
            9'd344: begin
                w_re = 10'sd13;
                w_im = -10'sd127;
            end
            9'd345: begin
                w_re = 10'sd5;
                w_im = -10'sd128;
            end
            9'd346: begin
                w_re = -10'sd3;
                w_im = -10'sd128;
            end
            9'd347: begin
                w_re = -10'sd11;
                w_im = -10'sd128;
            end
            9'd348: begin
                w_re = -10'sd19;
                w_im = -10'sd127;
            end
            9'd349: begin
                w_re = -10'sd27;
                w_im = -10'sd125;
            end
            9'd350: begin
                w_re = -10'sd34;
                w_im = -10'sd123;
            end
            9'd351: begin
                w_re = -10'sd42;
                w_im = -10'sd121;
            end
            9'd352: begin
                w_re = -10'sd49;
                w_im = -10'sd118;
            end
            9'd353: begin
                w_re = -10'sd56;
                w_im = -10'sd115;
            end
            9'd354: begin
                w_re = -10'sd63;
                w_im = -10'sd111;
            end
            9'd355: begin
                w_re = -10'sd70;
                w_im = -10'sd107;
            end
            9'd356: begin
                w_re = -10'sd76;
                w_im = -10'sd103;
            end
            9'd357: begin
                w_re = -10'sd82;
                w_im = -10'sd98;
            end
            9'd358: begin
                w_re = -10'sd88;
                w_im = -10'sd93;
            end
            9'd359: begin
                w_re = -10'sd94;
                w_im = -10'sd87;
            end
            9'd360: begin
                w_re = -10'sd99;
                w_im = -10'sd81;
            end
            9'd361: begin
                w_re = -10'sd104;
                w_im = -10'sd75;
            end
            9'd362: begin
                w_re = -10'sd108;
                w_im = -10'sd68;
            end
            9'd363: begin
                w_re = -10'sd112;
                w_im = -10'sd62;
            end
            9'd364: begin
                w_re = -10'sd116;
                w_im = -10'sd55;
            end
            9'd365: begin
                w_re = -10'sd119;
                w_im = -10'sd48;
            end
            9'd366: begin
                w_re = -10'sd122;
                w_im = -10'sd40;
            end
            9'd367: begin
                w_re = -10'sd124;
                w_im = -10'sd33;
            end
            9'd368: begin
                w_re = -10'sd126;
                w_im = -10'sd25;
            end
            9'd369: begin
                w_re = -10'sd127;
                w_im = -10'sd17;
            end
            9'd370: begin
                w_re = -10'sd128;
                w_im = -10'sd9;
            end
            9'd371: begin
                w_re = -10'sd128;
                w_im = -10'sd2;
            end
            9'd372: begin
                w_re = -10'sd128;
                w_im = 10'sd6;
            end
            9'd373: begin
                w_re = -10'sd127;
                w_im = 10'sd14;
            end
            9'd374: begin
                w_re = -10'sd126;
                w_im = 10'sd22;
            end
            9'd375: begin
                w_re = -10'sd125;
                w_im = 10'sd30;
            end
            9'd376: begin
                w_re = -10'sd122;
                w_im = 10'sd37;
            end
            9'd377: begin
                w_re = -10'sd120;
                w_im = 10'sd45;
            end
            9'd378: begin
                w_re = -10'sd117;
                w_im = 10'sd52;
            end
            9'd379: begin
                w_re = -10'sd114;
                w_im = 10'sd59;
            end
            9'd380: begin
                w_re = -10'sd110;
                w_im = 10'sd66;
            end
            9'd381: begin
                w_re = -10'sd106;
                w_im = 10'sd72;
            end
            9'd382: begin
                w_re = -10'sd101;
                w_im = 10'sd79;
            end
            9'd383: begin
                w_re = -10'sd96;
                w_im = 10'sd85;
            end
            9'd384: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd385: begin
                w_re = 10'sd128;
                w_im = -10'sd5;
            end
            9'd386: begin
                w_re = 10'sd128;
                w_im = -10'sd9;
            end
            9'd387: begin
                w_re = 10'sd127;
                w_im = -10'sd14;
            end
            9'd388: begin
                w_re = 10'sd127;
                w_im = -10'sd19;
            end
            9'd389: begin
                w_re = 10'sd126;
                w_im = -10'sd23;
            end
            9'd390: begin
                w_re = 10'sd125;
                w_im = -10'sd28;
            end
            9'd391: begin
                w_re = 10'sd124;
                w_im = -10'sd33;
            end
            9'd392: begin
                w_re = 10'sd122;
                w_im = -10'sd37;
            end
            9'd393: begin
                w_re = 10'sd121;
                w_im = -10'sd42;
            end
            9'd394: begin
                w_re = 10'sd119;
                w_im = -10'sd46;
            end
            9'd395: begin
                w_re = 10'sd118;
                w_im = -10'sd50;
            end
            9'd396: begin
                w_re = 10'sd116;
                w_im = -10'sd55;
            end
            9'd397: begin
                w_re = 10'sd114;
                w_im = -10'sd59;
            end
            9'd398: begin
                w_re = 10'sd111;
                w_im = -10'sd63;
            end
            9'd399: begin
                w_re = 10'sd109;
                w_im = -10'sd67;
            end
            9'd400: begin
                w_re = 10'sd106;
                w_im = -10'sd71;
            end
            9'd401: begin
                w_re = 10'sd104;
                w_im = -10'sd75;
            end
            9'd402: begin
                w_re = 10'sd101;
                w_im = -10'sd79;
            end
            9'd403: begin
                w_re = 10'sd98;
                w_im = -10'sd82;
            end
            9'd404: begin
                w_re = 10'sd95;
                w_im = -10'sd86;
            end
            9'd405: begin
                w_re = 10'sd92;
                w_im = -10'sd89;
            end
            9'd406: begin
                w_re = 10'sd88;
                w_im = -10'sd93;
            end
            9'd407: begin
                w_re = 10'sd85;
                w_im = -10'sd96;
            end
            9'd408: begin
                w_re = 10'sd81;
                w_im = -10'sd99;
            end
            9'd409: begin
                w_re = 10'sd78;
                w_im = -10'sd102;
            end
            9'd410: begin
                w_re = 10'sd74;
                w_im = -10'sd105;
            end
            9'd411: begin
                w_re = 10'sd70;
                w_im = -10'sd107;
            end
            9'd412: begin
                w_re = 10'sd66;
                w_im = -10'sd110;
            end
            9'd413: begin
                w_re = 10'sd62;
                w_im = -10'sd112;
            end
            9'd414: begin
                w_re = 10'sd58;
                w_im = -10'sd114;
            end
            9'd415: begin
                w_re = 10'sd53;
                w_im = -10'sd116;
            end
            9'd416: begin
                w_re = 10'sd49;
                w_im = -10'sd118;
            end
            9'd417: begin
                w_re = 10'sd45;
                w_im = -10'sd120;
            end
            9'd418: begin
                w_re = 10'sd40;
                w_im = -10'sd122;
            end
            9'd419: begin
                w_re = 10'sd36;
                w_im = -10'sd123;
            end
            9'd420: begin
                w_re = 10'sd31;
                w_im = -10'sd124;
            end
            9'd421: begin
                w_re = 10'sd27;
                w_im = -10'sd125;
            end
            9'd422: begin
                w_re = 10'sd22;
                w_im = -10'sd126;
            end
            9'd423: begin
                w_re = 10'sd17;
                w_im = -10'sd127;
            end
            9'd424: begin
                w_re = 10'sd13;
                w_im = -10'sd127;
            end
            9'd425: begin
                w_re = 10'sd8;
                w_im = -10'sd128;
            end
            9'd426: begin
                w_re = 10'sd3;
                w_im = -10'sd128;
            end
            9'd427: begin
                w_re = -10'sd2;
                w_im = -10'sd128;
            end
            9'd428: begin
                w_re = -10'sd6;
                w_im = -10'sd128;
            end
            9'd429: begin
                w_re = -10'sd11;
                w_im = -10'sd128;
            end
            9'd430: begin
                w_re = -10'sd16;
                w_im = -10'sd127;
            end
            9'd431: begin
                w_re = -10'sd20;
                w_im = -10'sd126;
            end
            9'd432: begin
                w_re = -10'sd25;
                w_im = -10'sd126;
            end
            9'd433: begin
                w_re = -10'sd30;
                w_im = -10'sd125;
            end
            9'd434: begin
                w_re = -10'sd34;
                w_im = -10'sd123;
            end
            9'd435: begin
                w_re = -10'sd39;
                w_im = -10'sd122;
            end
            9'd436: begin
                w_re = -10'sd43;
                w_im = -10'sd121;
            end
            9'd437: begin
                w_re = -10'sd48;
                w_im = -10'sd119;
            end
            9'd438: begin
                w_re = -10'sd52;
                w_im = -10'sd117;
            end
            9'd439: begin
                w_re = -10'sd56;
                w_im = -10'sd115;
            end
            9'd440: begin
                w_re = -10'sd60;
                w_im = -10'sd113;
            end
            9'd441: begin
                w_re = -10'sd64;
                w_im = -10'sd111;
            end
            9'd442: begin
                w_re = -10'sd68;
                w_im = -10'sd108;
            end
            9'd443: begin
                w_re = -10'sd72;
                w_im = -10'sd106;
            end
            9'd444: begin
                w_re = -10'sd76;
                w_im = -10'sd103;
            end
            9'd445: begin
                w_re = -10'sd80;
                w_im = -10'sd100;
            end
            9'd446: begin
                w_re = -10'sd84;
                w_im = -10'sd97;
            end
            9'd447: begin
                w_re = -10'sd87;
                w_im = -10'sd94;
            end
            9'd448: begin
                w_re = 10'sd128;
                w_im = 10'sd0;
            end
            9'd449: begin
                w_re = 10'sd128;
                w_im = -10'sd11;
            end
            9'd450: begin
                w_re = 10'sd126;
                w_im = -10'sd22;
            end
            9'd451: begin
                w_re = 10'sd124;
                w_im = -10'sd33;
            end
            9'd452: begin
                w_re = 10'sd121;
                w_im = -10'sd43;
            end
            9'd453: begin
                w_re = 10'sd116;
                w_im = -10'sd53;
            end
            9'd454: begin
                w_re = 10'sd111;
                w_im = -10'sd63;
            end
            9'd455: begin
                w_re = 10'sd106;
                w_im = -10'sd72;
            end
            9'd456: begin
                w_re = 10'sd99;
                w_im = -10'sd81;
            end
            9'd457: begin
                w_re = 10'sd92;
                w_im = -10'sd89;
            end
            9'd458: begin
                w_re = 10'sd84;
                w_im = -10'sd97;
            end
            9'd459: begin
                w_re = 10'sd75;
                w_im = -10'sd104;
            end
            9'd460: begin
                w_re = 10'sd66;
                w_im = -10'sd110;
            end
            9'd461: begin
                w_re = 10'sd56;
                w_im = -10'sd115;
            end
            9'd462: begin
                w_re = 10'sd46;
                w_im = -10'sd119;
            end
            9'd463: begin
                w_re = 10'sd36;
                w_im = -10'sd123;
            end
            9'd464: begin
                w_re = 10'sd25;
                w_im = -10'sd126;
            end
            9'd465: begin
                w_re = 10'sd14;
                w_im = -10'sd127;
            end
            9'd466: begin
                w_re = 10'sd3;
                w_im = -10'sd128;
            end
            9'd467: begin
                w_re = -10'sd8;
                w_im = -10'sd128;
            end
            9'd468: begin
                w_re = -10'sd19;
                w_im = -10'sd127;
            end
            9'd469: begin
                w_re = -10'sd30;
                w_im = -10'sd125;
            end
            9'd470: begin
                w_re = -10'sd40;
                w_im = -10'sd122;
            end
            9'd471: begin
                w_re = -10'sd50;
                w_im = -10'sd118;
            end
            9'd472: begin
                w_re = -10'sd60;
                w_im = -10'sd113;
            end
            9'd473: begin
                w_re = -10'sd70;
                w_im = -10'sd107;
            end
            9'd474: begin
                w_re = -10'sd79;
                w_im = -10'sd101;
            end
            9'd475: begin
                w_re = -10'sd87;
                w_im = -10'sd94;
            end
            9'd476: begin
                w_re = -10'sd95;
                w_im = -10'sd86;
            end
            9'd477: begin
                w_re = -10'sd102;
                w_im = -10'sd78;
            end
            9'd478: begin
                w_re = -10'sd108;
                w_im = -10'sd68;
            end
            9'd479: begin
                w_re = -10'sd114;
                w_im = -10'sd59;
            end
            9'd480: begin
                w_re = -10'sd118;
                w_im = -10'sd49;
            end
            9'd481: begin
                w_re = -10'sd122;
                w_im = -10'sd39;
            end
            9'd482: begin
                w_re = -10'sd125;
                w_im = -10'sd28;
            end
            9'd483: begin
                w_re = -10'sd127;
                w_im = -10'sd17;
            end
            9'd484: begin
                w_re = -10'sd128;
                w_im = -10'sd6;
            end
            9'd485: begin
                w_re = -10'sd128;
                w_im = 10'sd5;
            end
            9'd486: begin
                w_re = -10'sd127;
                w_im = 10'sd16;
            end
            9'd487: begin
                w_re = -10'sd125;
                w_im = 10'sd27;
            end
            9'd488: begin
                w_re = -10'sd122;
                w_im = 10'sd37;
            end
            9'd489: begin
                w_re = -10'sd119;
                w_im = 10'sd48;
            end
            9'd490: begin
                w_re = -10'sd114;
                w_im = 10'sd58;
            end
            9'd491: begin
                w_re = -10'sd109;
                w_im = 10'sd67;
            end
            9'd492: begin
                w_re = -10'sd103;
                w_im = 10'sd76;
            end
            9'd493: begin
                w_re = -10'sd96;
                w_im = 10'sd85;
            end
            9'd494: begin
                w_re = -10'sd88;
                w_im = 10'sd93;
            end
            9'd495: begin
                w_re = -10'sd80;
                w_im = 10'sd100;
            end
            9'd496: begin
                w_re = -10'sd71;
                w_im = 10'sd106;
            end
            9'd497: begin
                w_re = -10'sd62;
                w_im = 10'sd112;
            end
            9'd498: begin
                w_re = -10'sd52;
                w_im = 10'sd117;
            end
            9'd499: begin
                w_re = -10'sd42;
                w_im = 10'sd121;
            end
            9'd500: begin
                w_re = -10'sd31;
                w_im = 10'sd124;
            end
            9'd501: begin
                w_re = -10'sd20;
                w_im = 10'sd126;
            end
            9'd502: begin
                w_re = -10'sd9;
                w_im = 10'sd128;
            end
            9'd503: begin
                w_re = 10'sd2;
                w_im = 10'sd128;
            end
            9'd504: begin
                w_re = 10'sd13;
                w_im = 10'sd127;
            end
            9'd505: begin
                w_re = 10'sd23;
                w_im = 10'sd126;
            end
            9'd506: begin
                w_re = 10'sd34;
                w_im = 10'sd123;
            end
            9'd507: begin
                w_re = 10'sd45;
                w_im = 10'sd120;
            end
            9'd508: begin
                w_re = 10'sd55;
                w_im = 10'sd116;
            end
            9'd509: begin
                w_re = 10'sd64;
                w_im = 10'sd111;
            end
            9'd510: begin
                w_re = 10'sd74;
                w_im = 10'sd105;
            end
            9'd511: begin
                w_re = 10'sd82;
                w_im = 10'sd98;
            end

            // synopsys translate_off
            default: begin
                w_re = 10'sd0;
                w_im = 10'sd0;
            end
            // synopsys translate_on

        endcase
    end
endmodule
