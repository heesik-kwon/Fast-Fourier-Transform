`timescale 1ns / 1ps

module reverse #(
    parameter int N = 512,
    parameter int WIDTH = 13
) (
    input  logic signed [WIDTH-1:0] re_bfly22 [0:N-1],
    input  logic signed [WIDTH-1:0] im_bfly22 [0:N-1],
    output logic signed [WIDTH-1:0] re_dout[0:N-1],
    output logic signed [WIDTH-1:0] im_dout[0:N-1]
);

    // 비트 리버스 테이블
    localparam [8:0] bit_reverse_table [0:511] = '{
        9'd0,   9'd256, 9'd128, 9'd384, 9'd64,  9'd320, 9'd192, 9'd448,
        9'd32,  9'd288, 9'd160, 9'd416, 9'd96,  9'd352, 9'd224, 9'd480,
        9'd16,  9'd272, 9'd144, 9'd400, 9'd80,  9'd336, 9'd208, 9'd464,
        9'd48,  9'd304, 9'd176, 9'd432, 9'd112, 9'd368, 9'd240, 9'd496,
        9'd8,   9'd264, 9'd136, 9'd392, 9'd72,  9'd328, 9'd200, 9'd456,
        9'd40,  9'd296, 9'd168, 9'd424, 9'd104, 9'd360, 9'd232, 9'd488,
        9'd24,  9'd280, 9'd152, 9'd408, 9'd88,  9'd344, 9'd216, 9'd472,
        9'd56,  9'd312, 9'd184, 9'd440, 9'd120, 9'd376, 9'd248, 9'd504,
        9'd4,   9'd260, 9'd132, 9'd388, 9'd68,  9'd324, 9'd196, 9'd452,
        9'd36,  9'd292, 9'd164, 9'd420, 9'd100, 9'd356, 9'd228, 9'd484,
        9'd20,  9'd276, 9'd148, 9'd404, 9'd84,  9'd340, 9'd212, 9'd468,
        9'd52,  9'd308, 9'd180, 9'd436, 9'd116, 9'd372, 9'd244, 9'd500,
        9'd12,  9'd268, 9'd140, 9'd396, 9'd76,  9'd332, 9'd204, 9'd460,
        9'd44,  9'd300, 9'd172, 9'd428, 9'd108, 9'd364, 9'd236, 9'd492,
        9'd28,  9'd284, 9'd156, 9'd412, 9'd92,  9'd348, 9'd220, 9'd476,
        9'd60,  9'd316, 9'd188, 9'd444, 9'd124, 9'd380, 9'd252, 9'd508,
        9'd2,   9'd258, 9'd130, 9'd386, 9'd66,  9'd322, 9'd194, 9'd450,
        9'd34,  9'd290, 9'd162, 9'd418, 9'd98,  9'd354, 9'd226, 9'd482,
        9'd18,  9'd274, 9'd146, 9'd402, 9'd82,  9'd338, 9'd210, 9'd466,
        9'd50,  9'd306, 9'd178, 9'd434, 9'd114, 9'd370, 9'd242, 9'd498,
        9'd10,  9'd266, 9'd138, 9'd394, 9'd74,  9'd330, 9'd202, 9'd458,
        9'd42,  9'd298, 9'd170, 9'd426, 9'd106, 9'd362, 9'd234, 9'd490,
        9'd26,  9'd282, 9'd154, 9'd410, 9'd90,  9'd346, 9'd218, 9'd474,
        9'd58,  9'd314, 9'd186, 9'd442, 9'd122, 9'd378, 9'd250, 9'd506,
        9'd6,   9'd262, 9'd134, 9'd390, 9'd70,  9'd326, 9'd198, 9'd454,
        9'd38,  9'd294, 9'd166, 9'd422, 9'd102, 9'd358, 9'd230, 9'd486,
        9'd22,  9'd278, 9'd150, 9'd406, 9'd86,  9'd342, 9'd214, 9'd470,
        9'd54,  9'd310, 9'd182, 9'd438, 9'd118, 9'd374, 9'd246, 9'd502,
        9'd14,  9'd270, 9'd142, 9'd398, 9'd78,  9'd334, 9'd206, 9'd462,
        9'd46,  9'd302, 9'd174, 9'd430, 9'd110, 9'd366, 9'd238, 9'd494,
        9'd30,  9'd286, 9'd158, 9'd414, 9'd94,  9'd350, 9'd222, 9'd478,
        9'd62,  9'd318, 9'd190, 9'd446, 9'd126, 9'd382, 9'd254, 9'd510,
        9'd1,   9'd257, 9'd129, 9'd385, 9'd65,  9'd321, 9'd193, 9'd449,
        9'd33,  9'd289, 9'd161, 9'd417, 9'd97,  9'd353, 9'd225, 9'd481,
        9'd17,  9'd273, 9'd145, 9'd401, 9'd81,  9'd337, 9'd209, 9'd465,
        9'd49,  9'd305, 9'd177, 9'd433, 9'd113, 9'd369, 9'd241, 9'd497,
        9'd9,   9'd265, 9'd137, 9'd393, 9'd73,  9'd329, 9'd201, 9'd457,
        9'd41,  9'd297, 9'd169, 9'd425, 9'd105, 9'd361, 9'd233, 9'd489,
        9'd25,  9'd281, 9'd153, 9'd409, 9'd89,  9'd345, 9'd217, 9'd473,
        9'd57,  9'd313, 9'd185, 9'd441, 9'd121, 9'd377, 9'd249, 9'd505,
        9'd5,   9'd261, 9'd133, 9'd389, 9'd69,  9'd325, 9'd197, 9'd453,
        9'd37,  9'd293, 9'd165, 9'd421, 9'd101, 9'd357, 9'd229, 9'd485,
        9'd21,  9'd277, 9'd149, 9'd405, 9'd85,  9'd341, 9'd213, 9'd469,
        9'd53,  9'd309, 9'd181, 9'd437, 9'd117, 9'd373, 9'd245, 9'd501,
        9'd13,  9'd269, 9'd141, 9'd397, 9'd77,  9'd333, 9'd205, 9'd461,
        9'd45,  9'd301, 9'd173, 9'd429, 9'd109, 9'd365, 9'd237, 9'd493,
        9'd29,  9'd285, 9'd157, 9'd413, 9'd93,  9'd349, 9'd221, 9'd477,
        9'd61,  9'd317, 9'd189, 9'd445, 9'd125, 9'd381, 9'd253, 9'd509,
        9'd3,   9'd259, 9'd131, 9'd387, 9'd67,  9'd323, 9'd195, 9'd451,
        9'd35,  9'd291, 9'd163, 9'd419, 9'd99,  9'd355, 9'd227, 9'd483,
        9'd19,  9'd275, 9'd147, 9'd403, 9'd83,  9'd339, 9'd211, 9'd467,
        9'd51,  9'd307, 9'd179, 9'd435, 9'd115, 9'd371, 9'd243, 9'd499,
        9'd11,  9'd267, 9'd139, 9'd395, 9'd75,  9'd331, 9'd203, 9'd459,
        9'd43,  9'd299, 9'd171, 9'd427, 9'd107, 9'd363, 9'd235, 9'd491,
        9'd27,  9'd283, 9'd155, 9'd411, 9'd91,  9'd347, 9'd219, 9'd475,
        9'd59,  9'd315, 9'd187, 9'd443, 9'd123, 9'd379, 9'd251, 9'd507,
        9'd7,   9'd263, 9'd135, 9'd391, 9'd71,  9'd327, 9'd199, 9'd455,
        9'd39,  9'd295, 9'd167, 9'd423, 9'd103, 9'd359, 9'd231, 9'd487,
        9'd23,  9'd279, 9'd151, 9'd407, 9'd87,  9'd343, 9'd215, 9'd471,
        9'd55,  9'd311, 9'd183, 9'd439, 9'd119, 9'd375, 9'd247, 9'd503,
        9'd15,  9'd271, 9'd143, 9'd399, 9'd79,  9'd335, 9'd207, 9'd463,
        9'd47,  9'd303, 9'd175, 9'd431, 9'd111, 9'd367, 9'd239, 9'd495,
        9'd31,  9'd287, 9'd159, 9'd415, 9'd95,  9'd351, 9'd223, 9'd479,
        9'd63,  9'd319, 9'd191, 9'd447, 9'd127, 9'd383, 9'd255, 9'd511
    };

    genvar i;
    generate
        for (i = 0; i < N; i++) begin : GEN_ASSIGN
            assign re_dout[bit_reverse_table[i]] = re_bfly22[i];
            assign im_dout[bit_reverse_table[i]] = im_bfly22[i];
        end
    endgenerate

endmodule
